module controlunit(output regdst.
output jump,
output branch,
output memrd,
output memwr,
output aluop,
output memtoreg,
output regwr,
output alu8,
input [5:0] opcode
);





endmodule