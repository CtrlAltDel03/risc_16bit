module or32(
    output [31:0] out,
    input [31:0] a,b
);
assign {out}=a|b;

endmodule